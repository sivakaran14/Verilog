module bufif1gate(Y,A,B);
input A,B;
output Y;
bufif1 d1(Y,A,B);
endmodule
