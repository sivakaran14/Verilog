module tb_fulladder;
reg a,b,c;
wire s,d;
fulladder f1(.A(a),.B(b),.C(c),.S(s),.D(d));
initial 
begin         
a=1'b0;b=1'b0;c=1'b0;
#10 a=1'b0; b=1'b0;c=1'b1;
#10 a=1'b0; b=1'b1;c=1'b0;

#10 a=1'b0; b=1'b1;c=1'b1;
#10 a=1'b1; b=1'b0;c=1'b0;
#10 a=1'b1; b=1'b0;c=1'b1;
#10 a=1'b1; b=1'b1;c=1'b0;
#10 a=1'b1; b=1'b1;c=1'b1;
#100;$finish;
end
initial
begin
$dumpfile("tb_fulladder.vcd");
$dumpvars(0,tb_fulladder);
end
endmodule
