module bufgate(y,a);
input a;
output y;
buf b1(y,a);
endmodule
